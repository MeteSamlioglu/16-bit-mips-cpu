library verilog;
use verilog.vl_types.all;
entity test_registers is
end test_registers;
