library verilog;
use verilog.vl_types.all;
entity test_Mips is
end test_Mips;
