library verilog;
use verilog.vl_types.all;
entity test_instruction_memory is
end test_instruction_memory;
