library verilog;
use verilog.vl_types.all;
entity Alu_control_test is
end Alu_control_test;
