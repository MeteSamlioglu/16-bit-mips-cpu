library verilog;
use verilog.vl_types.all;
entity control_unit_test is
end control_unit_test;
