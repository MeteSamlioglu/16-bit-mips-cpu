library verilog;
use verilog.vl_types.all;
entity test_alu16bit is
end test_alu16bit;
